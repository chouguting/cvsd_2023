// list all paths to your design files
`include "../01_RTL/IOTDF.v"
`include "../01_RTL/inputReceiver.v"
`include "../01_RTL/desModule.v"
`include "../01_RTL/desKeyScheduler.v"
`include "../01_RTL/desFfunction.v"
`include "../01_RTL/outputModule.v"
`include "../01_RTL/crcModule.v"
`include "../01_RTL/binaryGrayConverter.v"

