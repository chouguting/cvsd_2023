module fisr ( // 4 dimensional vector dot product
    i_square_sum_u,  //
    o_isr,           // 1.11, unsign
    o_isr_shift_amt, // 
    o_isr_shift_dir
);
parameter S1_11_WIDTH = 13;
parameter S3_11_WIDTH = 15;
parameter S6_11_WIDTH = 18;

// parameter I_VEC_IM_WIDTH     = S1_11_WIDTH;
parameter SQUARE_SUM_WIDTH   = S6_11_WIDTH;
parameter SQUARE_SUM_U_WIDTH = SQUARE_SUM_WIDTH - 1;

// IO description
// input                          i_clk;
// input                          i_rst;

input  [SQUARE_SUM_U_WIDTH-1 : 0] i_square_sum_u;
output [S1_11_WIDTH-2        : 0] o_isr;
output [3 : 0]                    o_isr_shift_amt;
output                            o_isr_shift_dir;


// 17 bits, format: 6.11

// Instance of DW_lzd
// i_square_sum_u = [  00 00 00 . 00 | 00 00 00 00 | x ] ( if all 0's, last bit must be 1, underflow saturation)
//                [ 16                             0 ]

wire L1  = |i_square_sum_u[16 : 9];
wire R1  = |i_square_sum_u[8 : 1];
wire L1L = |i_square_sum_u[16 : 13];
wire R1L = |i_square_sum_u[8 : 5];
wire P1  = |i_square_sum_u[16 : 15]; 
wire P3  = |i_square_sum_u[12 : 11]; 
wire P5  = |i_square_sum_u[8 : 7]; 
wire P7  = |i_square_sum_u[4 : 3]; 

// wire L1R = |i_square_sum_u[12 : 9];
// wire R1R = |i_square_sum_u[4 : 1];
// wire P2 = |i_square_sum_u[14 : 13]; 
// wire P4 = |i_square_sum_u[10 : 9]; 
// wire P6 = |i_square_sum_u[6 : 5]; 
// wire P8 = |i_square_sum_u[2 : 1]; 

parameter RIGHT = 1'b0;
parameter LEFT  = 1'b1;
reg [4:0] shift_amt;
reg shift_dir;

always @(*) begin
    if(L1)begin
        if(L1L)begin
            if(P1)begin
                shift_amt = 5'd6;
                shift_dir = RIGHT;
            end
            else begin // P2
                shift_amt = 5'd4;
                shift_dir = RIGHT;
            end
        end
        else begin // L1R
            if(P3)begin
                shift_amt = 5'd2;
                shift_dir = RIGHT;
            end
            else begin // P4
                shift_amt = 5'd0;
                shift_dir = RIGHT;
            end
        end
    end
    else if(R1)begin
        if(R1L)begin
            if(P5)begin
                shift_amt = 5'd2;
                shift_dir = LEFT;
            end
            else begin // P6
                shift_amt = 5'd4;
                shift_dir = LEFT;
            end
        end
        else begin // R1R
            if(P7)begin
                shift_amt = 5'd6;
                shift_dir = LEFT;
            end
            else begin // P8
                shift_amt = 5'd8;
                shift_dir = LEFT;
            end
        end
    end 
    else begin
        shift_amt = 10;
        shift_dir = LEFT;
    end
end

// 0.1xxx or 0.x1xx format
// 17 bits, format: 6.11
wire [SQUARE_SUM_U_WIDTH-1 : 0] square_sum_u_shifted = (shift_dir == RIGHT) ? i_square_sum_u >> shift_amt : i_square_sum_u << shift_amt;

parameter a_width = 10; // format: .10 (fraction only)
wire [a_width-1 : 0] a = (~|i_square_sum_u)? {1'b1, 9'b0} : square_sum_u_shifted[SQUARE_SUM_U_WIDTH-1 -6 -: a_width]; // inverse square root input

// LUT 
wire [9:0] isr_frac [256:1023];
    assign isr_frac[256] = 10'b1111111111;
    assign isr_frac[257] = 10'b1111111100;
    assign isr_frac[258] = 10'b1111111000;
    assign isr_frac[259] = 10'b1111110100;
    assign isr_frac[260] = 10'b1111110000;
    assign isr_frac[261] = 10'b1111101100;
    assign isr_frac[262] = 10'b1111101000;
    assign isr_frac[263] = 10'b1111100100;
    assign isr_frac[264] = 10'b1111100000;
    assign isr_frac[265] = 10'b1111011100;
    assign isr_frac[266] = 10'b1111011001;
    assign isr_frac[267] = 10'b1111010101;
    assign isr_frac[268] = 10'b1111010001;
    assign isr_frac[269] = 10'b1111001101;
    assign isr_frac[270] = 10'b1111001010;
    assign isr_frac[271] = 10'b1111000110;
    assign isr_frac[272] = 10'b1111000010;
    assign isr_frac[273] = 10'b1110111111;
    assign isr_frac[274] = 10'b1110111011;
    assign isr_frac[275] = 10'b1110110111;
    assign isr_frac[276] = 10'b1110110100;
    assign isr_frac[277] = 10'b1110110000;
    assign isr_frac[278] = 10'b1110101101;
    assign isr_frac[279] = 10'b1110101001;
    assign isr_frac[280] = 10'b1110100110;
    assign isr_frac[281] = 10'b1110100010;
    assign isr_frac[282] = 10'b1110011111;
    assign isr_frac[283] = 10'b1110011011;
    assign isr_frac[284] = 10'b1110011000;
    assign isr_frac[285] = 10'b1110010101;
    assign isr_frac[286] = 10'b1110010001;
    assign isr_frac[287] = 10'b1110001110;
    assign isr_frac[288] = 10'b1110001010;
    assign isr_frac[289] = 10'b1110000111;
    assign isr_frac[290] = 10'b1110000100;
    assign isr_frac[291] = 10'b1110000000;
    assign isr_frac[292] = 10'b1101111101;
    assign isr_frac[293] = 10'b1101111010;
    assign isr_frac[294] = 10'b1101110111;
    assign isr_frac[295] = 10'b1101110011;
    assign isr_frac[296] = 10'b1101110000;
    assign isr_frac[297] = 10'b1101101101;
    assign isr_frac[298] = 10'b1101101010;
    assign isr_frac[299] = 10'b1101100111;
    assign isr_frac[300] = 10'b1101100011;
    assign isr_frac[301] = 10'b1101100000;
    assign isr_frac[302] = 10'b1101011101;
    assign isr_frac[303] = 10'b1101011010;
    assign isr_frac[304] = 10'b1101010111;
    assign isr_frac[305] = 10'b1101010100;
    assign isr_frac[306] = 10'b1101010001;
    assign isr_frac[307] = 10'b1101001110;
    assign isr_frac[308] = 10'b1101001011;
    assign isr_frac[309] = 10'b1101001000;
    assign isr_frac[310] = 10'b1101000101;
    assign isr_frac[311] = 10'b1101000010;
    assign isr_frac[312] = 10'b1100111111;
    assign isr_frac[313] = 10'b1100111100;
    assign isr_frac[314] = 10'b1100111001;
    assign isr_frac[315] = 10'b1100110110;
    assign isr_frac[316] = 10'b1100110011;
    assign isr_frac[317] = 10'b1100110000;
    assign isr_frac[318] = 10'b1100101101;
    assign isr_frac[319] = 10'b1100101010;
    assign isr_frac[320] = 10'b1100100111;
    assign isr_frac[321] = 10'b1100100100;
    assign isr_frac[322] = 10'b1100100010;
    assign isr_frac[323] = 10'b1100011111;
    assign isr_frac[324] = 10'b1100011100;
    assign isr_frac[325] = 10'b1100011001;
    assign isr_frac[326] = 10'b1100010110;
    assign isr_frac[327] = 10'b1100010100;
    assign isr_frac[328] = 10'b1100010001;
    assign isr_frac[329] = 10'b1100001110;
    assign isr_frac[330] = 10'b1100001011;
    assign isr_frac[331] = 10'b1100001001;
    assign isr_frac[332] = 10'b1100000110;
    assign isr_frac[333] = 10'b1100000011;
    assign isr_frac[334] = 10'b1100000000;
    assign isr_frac[335] = 10'b1011111110;
    assign isr_frac[336] = 10'b1011111011;
    assign isr_frac[337] = 10'b1011111000;
    assign isr_frac[338] = 10'b1011110110;
    assign isr_frac[339] = 10'b1011110011;
    assign isr_frac[340] = 10'b1011110001;
    assign isr_frac[341] = 10'b1011101110;
    assign isr_frac[342] = 10'b1011101011;
    assign isr_frac[343] = 10'b1011101001;
    assign isr_frac[344] = 10'b1011100110;
    assign isr_frac[345] = 10'b1011100100;
    assign isr_frac[346] = 10'b1011100001;
    assign isr_frac[347] = 10'b1011011111;
    assign isr_frac[348] = 10'b1011011100;
    assign isr_frac[349] = 10'b1011011010;
    assign isr_frac[350] = 10'b1011010111;
    assign isr_frac[351] = 10'b1011010101;
    assign isr_frac[352] = 10'b1011010010;
    assign isr_frac[353] = 10'b1011010000;
    assign isr_frac[354] = 10'b1011001101;
    assign isr_frac[355] = 10'b1011001011;
    assign isr_frac[356] = 10'b1011001000;
    assign isr_frac[357] = 10'b1011000110;
    assign isr_frac[358] = 10'b1011000011;
    assign isr_frac[359] = 10'b1011000001;
    assign isr_frac[360] = 10'b1010111111;
    assign isr_frac[361] = 10'b1010111100;
    assign isr_frac[362] = 10'b1010111010;
    assign isr_frac[363] = 10'b1010110111;
    assign isr_frac[364] = 10'b1010110101;
    assign isr_frac[365] = 10'b1010110011;
    assign isr_frac[366] = 10'b1010110000;
    assign isr_frac[367] = 10'b1010101110;
    assign isr_frac[368] = 10'b1010101100;
    assign isr_frac[369] = 10'b1010101001;
    assign isr_frac[370] = 10'b1010100111;
    assign isr_frac[371] = 10'b1010100101;
    assign isr_frac[372] = 10'b1010100010;
    assign isr_frac[373] = 10'b1010100000;
    assign isr_frac[374] = 10'b1010011110;
    assign isr_frac[375] = 10'b1010011100;
    assign isr_frac[376] = 10'b1010011001;
    assign isr_frac[377] = 10'b1010010111;
    assign isr_frac[378] = 10'b1010010101;
    assign isr_frac[379] = 10'b1010010011;
    assign isr_frac[380] = 10'b1010010000;
    assign isr_frac[381] = 10'b1010001110;
    assign isr_frac[382] = 10'b1010001100;
    assign isr_frac[383] = 10'b1010001010;
    assign isr_frac[384] = 10'b1010001000;
    assign isr_frac[385] = 10'b1010000110;
    assign isr_frac[386] = 10'b1010000011;
    assign isr_frac[387] = 10'b1010000001;
    assign isr_frac[388] = 10'b1001111111;
    assign isr_frac[389] = 10'b1001111101;
    assign isr_frac[390] = 10'b1001111011;
    assign isr_frac[391] = 10'b1001111001;
    assign isr_frac[392] = 10'b1001110111;
    assign isr_frac[393] = 10'b1001110100;
    assign isr_frac[394] = 10'b1001110010;
    assign isr_frac[395] = 10'b1001110000;
    assign isr_frac[396] = 10'b1001101110;
    assign isr_frac[397] = 10'b1001101100;
    assign isr_frac[398] = 10'b1001101010;
    assign isr_frac[399] = 10'b1001101000;
    assign isr_frac[400] = 10'b1001100110;
    assign isr_frac[401] = 10'b1001100100;
    assign isr_frac[402] = 10'b1001100010;
    assign isr_frac[403] = 10'b1001100000;
    assign isr_frac[404] = 10'b1001011110;
    assign isr_frac[405] = 10'b1001011100;
    assign isr_frac[406] = 10'b1001011010;
    assign isr_frac[407] = 10'b1001011000;
    assign isr_frac[408] = 10'b1001010110;
    assign isr_frac[409] = 10'b1001010100;
    assign isr_frac[410] = 10'b1001010010;
    assign isr_frac[411] = 10'b1001010000;
    assign isr_frac[412] = 10'b1001001110;
    assign isr_frac[413] = 10'b1001001100;
    assign isr_frac[414] = 10'b1001001010;
    assign isr_frac[415] = 10'b1001001000;
    assign isr_frac[416] = 10'b1001000110;
    assign isr_frac[417] = 10'b1001000100;
    assign isr_frac[418] = 10'b1001000010;
    assign isr_frac[419] = 10'b1001000000;
    assign isr_frac[420] = 10'b1000111110;
    assign isr_frac[421] = 10'b1000111101;
    assign isr_frac[422] = 10'b1000111011;
    assign isr_frac[423] = 10'b1000111001;
    assign isr_frac[424] = 10'b1000110111;
    assign isr_frac[425] = 10'b1000110101;
    assign isr_frac[426] = 10'b1000110011;
    assign isr_frac[427] = 10'b1000110001;
    assign isr_frac[428] = 10'b1000101111;
    assign isr_frac[429] = 10'b1000101110;
    assign isr_frac[430] = 10'b1000101100;
    assign isr_frac[431] = 10'b1000101010;
    assign isr_frac[432] = 10'b1000101000;
    assign isr_frac[433] = 10'b1000100110;
    assign isr_frac[434] = 10'b1000100100;
    assign isr_frac[435] = 10'b1000100011;
    assign isr_frac[436] = 10'b1000100001;
    assign isr_frac[437] = 10'b1000011111;
    assign isr_frac[438] = 10'b1000011101;
    assign isr_frac[439] = 10'b1000011011;
    assign isr_frac[440] = 10'b1000011010;
    assign isr_frac[441] = 10'b1000011000;
    assign isr_frac[442] = 10'b1000010110;
    assign isr_frac[443] = 10'b1000010100;
    assign isr_frac[444] = 10'b1000010011;
    assign isr_frac[445] = 10'b1000010001;
    assign isr_frac[446] = 10'b1000001111;
    assign isr_frac[447] = 10'b1000001101;
    assign isr_frac[448] = 10'b1000001100;
    assign isr_frac[449] = 10'b1000001010;
    assign isr_frac[450] = 10'b1000001000;
    assign isr_frac[451] = 10'b1000000110;
    assign isr_frac[452] = 10'b1000000101;
    assign isr_frac[453] = 10'b1000000011;
    assign isr_frac[454] = 10'b1000000001;
    assign isr_frac[455] = 10'b1000000000;
    assign isr_frac[456] = 10'b0111111110;
    assign isr_frac[457] = 10'b0111111100;
    assign isr_frac[458] = 10'b0111111011;
    assign isr_frac[459] = 10'b0111111001;
    assign isr_frac[460] = 10'b0111110111;
    assign isr_frac[461] = 10'b0111110110;
    assign isr_frac[462] = 10'b0111110100;
    assign isr_frac[463] = 10'b0111110010;
    assign isr_frac[464] = 10'b0111110001;
    assign isr_frac[465] = 10'b0111101111;
    assign isr_frac[466] = 10'b0111101101;
    assign isr_frac[467] = 10'b0111101100;
    assign isr_frac[468] = 10'b0111101010;
    assign isr_frac[469] = 10'b0111101001;
    assign isr_frac[470] = 10'b0111100111;
    assign isr_frac[471] = 10'b0111100101;
    assign isr_frac[472] = 10'b0111100100;
    assign isr_frac[473] = 10'b0111100010;
    assign isr_frac[474] = 10'b0111100001;
    assign isr_frac[475] = 10'b0111011111;
    assign isr_frac[476] = 10'b0111011101;
    assign isr_frac[477] = 10'b0111011100;
    assign isr_frac[478] = 10'b0111011010;
    assign isr_frac[479] = 10'b0111011001;
    assign isr_frac[480] = 10'b0111010111;
    assign isr_frac[481] = 10'b0111010110;
    assign isr_frac[482] = 10'b0111010100;
    assign isr_frac[483] = 10'b0111010010;
    assign isr_frac[484] = 10'b0111010001;
    assign isr_frac[485] = 10'b0111001111;
    assign isr_frac[486] = 10'b0111001110;
    assign isr_frac[487] = 10'b0111001100;
    assign isr_frac[488] = 10'b0111001011;
    assign isr_frac[489] = 10'b0111001001;
    assign isr_frac[490] = 10'b0111001000;
    assign isr_frac[491] = 10'b0111000110;
    assign isr_frac[492] = 10'b0111000101;
    assign isr_frac[493] = 10'b0111000011;
    assign isr_frac[494] = 10'b0111000010;
    assign isr_frac[495] = 10'b0111000000;
    assign isr_frac[496] = 10'b0110111111;
    assign isr_frac[497] = 10'b0110111101;
    assign isr_frac[498] = 10'b0110111100;
    assign isr_frac[499] = 10'b0110111010;
    assign isr_frac[500] = 10'b0110111001;
    assign isr_frac[501] = 10'b0110110111;
    assign isr_frac[502] = 10'b0110110110;
    assign isr_frac[503] = 10'b0110110101;
    assign isr_frac[504] = 10'b0110110011;
    assign isr_frac[505] = 10'b0110110010;
    assign isr_frac[506] = 10'b0110110000;
    assign isr_frac[507] = 10'b0110101111;
    assign isr_frac[508] = 10'b0110101101;
    assign isr_frac[509] = 10'b0110101100;
    assign isr_frac[510] = 10'b0110101010;
    assign isr_frac[511] = 10'b0110101001;
    assign isr_frac[512] = 10'b0110101000;
    assign isr_frac[513] = 10'b0110100110;
    assign isr_frac[514] = 10'b0110100101;
    assign isr_frac[515] = 10'b0110100011;
    assign isr_frac[516] = 10'b0110100010;
    assign isr_frac[517] = 10'b0110100001;
    assign isr_frac[518] = 10'b0110011111;
    assign isr_frac[519] = 10'b0110011110;
    assign isr_frac[520] = 10'b0110011100;
    assign isr_frac[521] = 10'b0110011011;
    assign isr_frac[522] = 10'b0110011010;
    assign isr_frac[523] = 10'b0110011000;
    assign isr_frac[524] = 10'b0110010111;
    assign isr_frac[525] = 10'b0110010110;
    assign isr_frac[526] = 10'b0110010100;
    assign isr_frac[527] = 10'b0110010011;
    assign isr_frac[528] = 10'b0110010010;
    assign isr_frac[529] = 10'b0110010000;
    assign isr_frac[530] = 10'b0110001111;
    assign isr_frac[531] = 10'b0110001110;
    assign isr_frac[532] = 10'b0110001100;
    assign isr_frac[533] = 10'b0110001011;
    assign isr_frac[534] = 10'b0110001010;
    assign isr_frac[535] = 10'b0110001000;
    assign isr_frac[536] = 10'b0110000111;
    assign isr_frac[537] = 10'b0110000110;
    assign isr_frac[538] = 10'b0110000100;
    assign isr_frac[539] = 10'b0110000011;
    assign isr_frac[540] = 10'b0110000010;
    assign isr_frac[541] = 10'b0110000000;
    assign isr_frac[542] = 10'b0101111111;
    assign isr_frac[543] = 10'b0101111110;
    assign isr_frac[544] = 10'b0101111100;
    assign isr_frac[545] = 10'b0101111011;
    assign isr_frac[546] = 10'b0101111010;
    assign isr_frac[547] = 10'b0101111001;
    assign isr_frac[548] = 10'b0101110111;
    assign isr_frac[549] = 10'b0101110110;
    assign isr_frac[550] = 10'b0101110101;
    assign isr_frac[551] = 10'b0101110011;
    assign isr_frac[552] = 10'b0101110010;
    assign isr_frac[553] = 10'b0101110001;
    assign isr_frac[554] = 10'b0101110000;
    assign isr_frac[555] = 10'b0101101110;
    assign isr_frac[556] = 10'b0101101101;
    assign isr_frac[557] = 10'b0101101100;
    assign isr_frac[558] = 10'b0101101011;
    assign isr_frac[559] = 10'b0101101001;
    assign isr_frac[560] = 10'b0101101000;
    assign isr_frac[561] = 10'b0101100111;
    assign isr_frac[562] = 10'b0101100110;
    assign isr_frac[563] = 10'b0101100101;
    assign isr_frac[564] = 10'b0101100011;
    assign isr_frac[565] = 10'b0101100010;
    assign isr_frac[566] = 10'b0101100001;
    assign isr_frac[567] = 10'b0101100000;
    assign isr_frac[568] = 10'b0101011110;
    assign isr_frac[569] = 10'b0101011101;
    assign isr_frac[570] = 10'b0101011100;
    assign isr_frac[571] = 10'b0101011011;
    assign isr_frac[572] = 10'b0101011010;
    assign isr_frac[573] = 10'b0101011000;
    assign isr_frac[574] = 10'b0101010111;
    assign isr_frac[575] = 10'b0101010110;
    assign isr_frac[576] = 10'b0101010101;
    assign isr_frac[577] = 10'b0101010100;
    assign isr_frac[578] = 10'b0101010010;
    assign isr_frac[579] = 10'b0101010001;
    assign isr_frac[580] = 10'b0101010000;
    assign isr_frac[581] = 10'b0101001111;
    assign isr_frac[582] = 10'b0101001110;
    assign isr_frac[583] = 10'b0101001101;
    assign isr_frac[584] = 10'b0101001011;
    assign isr_frac[585] = 10'b0101001010;
    assign isr_frac[586] = 10'b0101001001;
    assign isr_frac[587] = 10'b0101001000;
    assign isr_frac[588] = 10'b0101000111;
    assign isr_frac[589] = 10'b0101000110;
    assign isr_frac[590] = 10'b0101000101;
    assign isr_frac[591] = 10'b0101000011;
    assign isr_frac[592] = 10'b0101000010;
    assign isr_frac[593] = 10'b0101000001;
    assign isr_frac[594] = 10'b0101000000;
    assign isr_frac[595] = 10'b0100111111;
    assign isr_frac[596] = 10'b0100111110;
    assign isr_frac[597] = 10'b0100111101;
    assign isr_frac[598] = 10'b0100111011;
    assign isr_frac[599] = 10'b0100111010;
    assign isr_frac[600] = 10'b0100111001;
    assign isr_frac[601] = 10'b0100111000;
    assign isr_frac[602] = 10'b0100110111;
    assign isr_frac[603] = 10'b0100110110;
    assign isr_frac[604] = 10'b0100110101;
    assign isr_frac[605] = 10'b0100110100;
    assign isr_frac[606] = 10'b0100110011;
    assign isr_frac[607] = 10'b0100110010;
    assign isr_frac[608] = 10'b0100110000;
    assign isr_frac[609] = 10'b0100101111;
    assign isr_frac[610] = 10'b0100101110;
    assign isr_frac[611] = 10'b0100101101;
    assign isr_frac[612] = 10'b0100101100;
    assign isr_frac[613] = 10'b0100101011;
    assign isr_frac[614] = 10'b0100101010;
    assign isr_frac[615] = 10'b0100101001;
    assign isr_frac[616] = 10'b0100101000;
    assign isr_frac[617] = 10'b0100100111;
    assign isr_frac[618] = 10'b0100100110;
    assign isr_frac[619] = 10'b0100100101;
    assign isr_frac[620] = 10'b0100100011;
    assign isr_frac[621] = 10'b0100100010;
    assign isr_frac[622] = 10'b0100100001;
    assign isr_frac[623] = 10'b0100100000;
    assign isr_frac[624] = 10'b0100011111;
    assign isr_frac[625] = 10'b0100011110;
    assign isr_frac[626] = 10'b0100011101;
    assign isr_frac[627] = 10'b0100011100;
    assign isr_frac[628] = 10'b0100011011;
    assign isr_frac[629] = 10'b0100011010;
    assign isr_frac[630] = 10'b0100011001;
    assign isr_frac[631] = 10'b0100011000;
    assign isr_frac[632] = 10'b0100010111;
    assign isr_frac[633] = 10'b0100010110;
    assign isr_frac[634] = 10'b0100010101;
    assign isr_frac[635] = 10'b0100010100;
    assign isr_frac[636] = 10'b0100010011;
    assign isr_frac[637] = 10'b0100010010;
    assign isr_frac[638] = 10'b0100010001;
    assign isr_frac[639] = 10'b0100010000;
    assign isr_frac[640] = 10'b0100001111;
    assign isr_frac[641] = 10'b0100001110;
    assign isr_frac[642] = 10'b0100001101;
    assign isr_frac[643] = 10'b0100001100;
    assign isr_frac[644] = 10'b0100001011;
    assign isr_frac[645] = 10'b0100001010;
    assign isr_frac[646] = 10'b0100001001;
    assign isr_frac[647] = 10'b0100001000;
    assign isr_frac[648] = 10'b0100000111;
    assign isr_frac[649] = 10'b0100000110;
    assign isr_frac[650] = 10'b0100000101;
    assign isr_frac[651] = 10'b0100000100;
    assign isr_frac[652] = 10'b0100000011;
    assign isr_frac[653] = 10'b0100000010;
    assign isr_frac[654] = 10'b0100000001;
    assign isr_frac[655] = 10'b0100000000;
    assign isr_frac[656] = 10'b0011111111;
    assign isr_frac[657] = 10'b0011111110;
    assign isr_frac[658] = 10'b0011111101;
    assign isr_frac[659] = 10'b0011111100;
    assign isr_frac[660] = 10'b0011111011;
    assign isr_frac[661] = 10'b0011111010;
    assign isr_frac[662] = 10'b0011111001;
    assign isr_frac[663] = 10'b0011111000;
    assign isr_frac[664] = 10'b0011110111;
    assign isr_frac[665] = 10'b0011110110;
    assign isr_frac[666] = 10'b0011110101;
    assign isr_frac[667] = 10'b0011110100;
    assign isr_frac[668] = 10'b0011110011;
    assign isr_frac[669] = 10'b0011110010;
    assign isr_frac[670] = 10'b0011110001;
    assign isr_frac[671] = 10'b0011110000;
    assign isr_frac[672] = 10'b0011110000;
    assign isr_frac[673] = 10'b0011101111;
    assign isr_frac[674] = 10'b0011101110;
    assign isr_frac[675] = 10'b0011101101;
    assign isr_frac[676] = 10'b0011101100;
    assign isr_frac[677] = 10'b0011101011;
    assign isr_frac[678] = 10'b0011101010;
    assign isr_frac[679] = 10'b0011101001;
    assign isr_frac[680] = 10'b0011101000;
    assign isr_frac[681] = 10'b0011100111;
    assign isr_frac[682] = 10'b0011100110;
    assign isr_frac[683] = 10'b0011100101;
    assign isr_frac[684] = 10'b0011100100;
    assign isr_frac[685] = 10'b0011100100;
    assign isr_frac[686] = 10'b0011100011;
    assign isr_frac[687] = 10'b0011100010;
    assign isr_frac[688] = 10'b0011100001;
    assign isr_frac[689] = 10'b0011100000;
    assign isr_frac[690] = 10'b0011011111;
    assign isr_frac[691] = 10'b0011011110;
    assign isr_frac[692] = 10'b0011011101;
    assign isr_frac[693] = 10'b0011011100;
    assign isr_frac[694] = 10'b0011011011;
    assign isr_frac[695] = 10'b0011011010;
    assign isr_frac[696] = 10'b0011011010;
    assign isr_frac[697] = 10'b0011011001;
    assign isr_frac[698] = 10'b0011011000;
    assign isr_frac[699] = 10'b0011010111;
    assign isr_frac[700] = 10'b0011010110;
    assign isr_frac[701] = 10'b0011010101;
    assign isr_frac[702] = 10'b0011010100;
    assign isr_frac[703] = 10'b0011010011;
    assign isr_frac[704] = 10'b0011010010;
    assign isr_frac[705] = 10'b0011010010;
    assign isr_frac[706] = 10'b0011010001;
    assign isr_frac[707] = 10'b0011010000;
    assign isr_frac[708] = 10'b0011001111;
    assign isr_frac[709] = 10'b0011001110;
    assign isr_frac[710] = 10'b0011001101;
    assign isr_frac[711] = 10'b0011001100;
    assign isr_frac[712] = 10'b0011001100;
    assign isr_frac[713] = 10'b0011001011;
    assign isr_frac[714] = 10'b0011001010;
    assign isr_frac[715] = 10'b0011001001;
    assign isr_frac[716] = 10'b0011001000;
    assign isr_frac[717] = 10'b0011000111;
    assign isr_frac[718] = 10'b0011000110;
    assign isr_frac[719] = 10'b0011000110;
    assign isr_frac[720] = 10'b0011000101;
    assign isr_frac[721] = 10'b0011000100;
    assign isr_frac[722] = 10'b0011000011;
    assign isr_frac[723] = 10'b0011000010;
    assign isr_frac[724] = 10'b0011000001;
    assign isr_frac[725] = 10'b0011000000;
    assign isr_frac[726] = 10'b0011000000;
    assign isr_frac[727] = 10'b0010111111;
    assign isr_frac[728] = 10'b0010111110;
    assign isr_frac[729] = 10'b0010111101;
    assign isr_frac[730] = 10'b0010111100;
    assign isr_frac[731] = 10'b0010111011;
    assign isr_frac[732] = 10'b0010111011;
    assign isr_frac[733] = 10'b0010111010;
    assign isr_frac[734] = 10'b0010111001;
    assign isr_frac[735] = 10'b0010111000;
    assign isr_frac[736] = 10'b0010110111;
    assign isr_frac[737] = 10'b0010110111;
    assign isr_frac[738] = 10'b0010110110;
    assign isr_frac[739] = 10'b0010110101;
    assign isr_frac[740] = 10'b0010110100;
    assign isr_frac[741] = 10'b0010110011;
    assign isr_frac[742] = 10'b0010110010;
    assign isr_frac[743] = 10'b0010110010;
    assign isr_frac[744] = 10'b0010110001;
    assign isr_frac[745] = 10'b0010110000;
    assign isr_frac[746] = 10'b0010101111;
    assign isr_frac[747] = 10'b0010101110;
    assign isr_frac[748] = 10'b0010101110;
    assign isr_frac[749] = 10'b0010101101;
    assign isr_frac[750] = 10'b0010101100;
    assign isr_frac[751] = 10'b0010101011;
    assign isr_frac[752] = 10'b0010101010;
    assign isr_frac[753] = 10'b0010101010;
    assign isr_frac[754] = 10'b0010101001;
    assign isr_frac[755] = 10'b0010101000;
    assign isr_frac[756] = 10'b0010100111;
    assign isr_frac[757] = 10'b0010100110;
    assign isr_frac[758] = 10'b0010100110;
    assign isr_frac[759] = 10'b0010100101;
    assign isr_frac[760] = 10'b0010100100;
    assign isr_frac[761] = 10'b0010100011;
    assign isr_frac[762] = 10'b0010100011;
    assign isr_frac[763] = 10'b0010100010;
    assign isr_frac[764] = 10'b0010100001;
    assign isr_frac[765] = 10'b0010100000;
    assign isr_frac[766] = 10'b0010011111;
    assign isr_frac[767] = 10'b0010011111;
    assign isr_frac[768] = 10'b0010011110;
    assign isr_frac[769] = 10'b0010011101;
    assign isr_frac[770] = 10'b0010011100;
    assign isr_frac[771] = 10'b0010011100;
    assign isr_frac[772] = 10'b0010011011;
    assign isr_frac[773] = 10'b0010011010;
    assign isr_frac[774] = 10'b0010011001;
    assign isr_frac[775] = 10'b0010011001;
    assign isr_frac[776] = 10'b0010011000;
    assign isr_frac[777] = 10'b0010010111;
    assign isr_frac[778] = 10'b0010010110;
    assign isr_frac[779] = 10'b0010010110;
    assign isr_frac[780] = 10'b0010010101;
    assign isr_frac[781] = 10'b0010010100;
    assign isr_frac[782] = 10'b0010010011;
    assign isr_frac[783] = 10'b0010010011;
    assign isr_frac[784] = 10'b0010010010;
    assign isr_frac[785] = 10'b0010010001;
    assign isr_frac[786] = 10'b0010010000;
    assign isr_frac[787] = 10'b0010010000;
    assign isr_frac[788] = 10'b0010001111;
    assign isr_frac[789] = 10'b0010001110;
    assign isr_frac[790] = 10'b0010001101;
    assign isr_frac[791] = 10'b0010001101;
    assign isr_frac[792] = 10'b0010001100;
    assign isr_frac[793] = 10'b0010001011;
    assign isr_frac[794] = 10'b0010001010;
    assign isr_frac[795] = 10'b0010001010;
    assign isr_frac[796] = 10'b0010001001;
    assign isr_frac[797] = 10'b0010001000;
    assign isr_frac[798] = 10'b0010000111;
    assign isr_frac[799] = 10'b0010000111;
    assign isr_frac[800] = 10'b0010000110;
    assign isr_frac[801] = 10'b0010000101;
    assign isr_frac[802] = 10'b0010000101;
    assign isr_frac[803] = 10'b0010000100;
    assign isr_frac[804] = 10'b0010000011;
    assign isr_frac[805] = 10'b0010000010;
    assign isr_frac[806] = 10'b0010000010;
    assign isr_frac[807] = 10'b0010000001;
    assign isr_frac[808] = 10'b0010000000;
    assign isr_frac[809] = 10'b0010000000;
    assign isr_frac[810] = 10'b0001111111;
    assign isr_frac[811] = 10'b0001111110;
    assign isr_frac[812] = 10'b0001111101;
    assign isr_frac[813] = 10'b0001111101;
    assign isr_frac[814] = 10'b0001111100;
    assign isr_frac[815] = 10'b0001111011;
    assign isr_frac[816] = 10'b0001111011;
    assign isr_frac[817] = 10'b0001111010;
    assign isr_frac[818] = 10'b0001111001;
    assign isr_frac[819] = 10'b0001111001;
    assign isr_frac[820] = 10'b0001111000;
    assign isr_frac[821] = 10'b0001110111;
    assign isr_frac[822] = 10'b0001110110;
    assign isr_frac[823] = 10'b0001110110;
    assign isr_frac[824] = 10'b0001110101;
    assign isr_frac[825] = 10'b0001110100;
    assign isr_frac[826] = 10'b0001110100;
    assign isr_frac[827] = 10'b0001110011;
    assign isr_frac[828] = 10'b0001110010;
    assign isr_frac[829] = 10'b0001110010;
    assign isr_frac[830] = 10'b0001110001;
    assign isr_frac[831] = 10'b0001110000;
    assign isr_frac[832] = 10'b0001110000;
    assign isr_frac[833] = 10'b0001101111;
    assign isr_frac[834] = 10'b0001101110;
    assign isr_frac[835] = 10'b0001101101;
    assign isr_frac[836] = 10'b0001101101;
    assign isr_frac[837] = 10'b0001101100;
    assign isr_frac[838] = 10'b0001101011;
    assign isr_frac[839] = 10'b0001101011;
    assign isr_frac[840] = 10'b0001101010;
    assign isr_frac[841] = 10'b0001101001;
    assign isr_frac[842] = 10'b0001101001;
    assign isr_frac[843] = 10'b0001101000;
    assign isr_frac[844] = 10'b0001100111;
    assign isr_frac[845] = 10'b0001100111;
    assign isr_frac[846] = 10'b0001100110;
    assign isr_frac[847] = 10'b0001100101;
    assign isr_frac[848] = 10'b0001100101;
    assign isr_frac[849] = 10'b0001100100;
    assign isr_frac[850] = 10'b0001100011;
    assign isr_frac[851] = 10'b0001100011;
    assign isr_frac[852] = 10'b0001100010;
    assign isr_frac[853] = 10'b0001100001;
    assign isr_frac[854] = 10'b0001100001;
    assign isr_frac[855] = 10'b0001100000;
    assign isr_frac[856] = 10'b0001011111;
    assign isr_frac[857] = 10'b0001011111;
    assign isr_frac[858] = 10'b0001011110;
    assign isr_frac[859] = 10'b0001011110;
    assign isr_frac[860] = 10'b0001011101;
    assign isr_frac[861] = 10'b0001011100;
    assign isr_frac[862] = 10'b0001011100;
    assign isr_frac[863] = 10'b0001011011;
    assign isr_frac[864] = 10'b0001011010;
    assign isr_frac[865] = 10'b0001011010;
    assign isr_frac[866] = 10'b0001011001;
    assign isr_frac[867] = 10'b0001011000;
    assign isr_frac[868] = 10'b0001011000;
    assign isr_frac[869] = 10'b0001010111;
    assign isr_frac[870] = 10'b0001010110;
    assign isr_frac[871] = 10'b0001010110;
    assign isr_frac[872] = 10'b0001010101;
    assign isr_frac[873] = 10'b0001010101;
    assign isr_frac[874] = 10'b0001010100;
    assign isr_frac[875] = 10'b0001010011;
    assign isr_frac[876] = 10'b0001010011;
    assign isr_frac[877] = 10'b0001010010;
    assign isr_frac[878] = 10'b0001010001;
    assign isr_frac[879] = 10'b0001010001;
    assign isr_frac[880] = 10'b0001010000;
    assign isr_frac[881] = 10'b0001001111;
    assign isr_frac[882] = 10'b0001001111;
    assign isr_frac[883] = 10'b0001001110;
    assign isr_frac[884] = 10'b0001001110;
    assign isr_frac[885] = 10'b0001001101;
    assign isr_frac[886] = 10'b0001001100;
    assign isr_frac[887] = 10'b0001001100;
    assign isr_frac[888] = 10'b0001001011;
    assign isr_frac[889] = 10'b0001001011;
    assign isr_frac[890] = 10'b0001001010;
    assign isr_frac[891] = 10'b0001001001;
    assign isr_frac[892] = 10'b0001001001;
    assign isr_frac[893] = 10'b0001001000;
    assign isr_frac[894] = 10'b0001000111;
    assign isr_frac[895] = 10'b0001000111;
    assign isr_frac[896] = 10'b0001000110;
    assign isr_frac[897] = 10'b0001000110;
    assign isr_frac[898] = 10'b0001000101;
    assign isr_frac[899] = 10'b0001000100;
    assign isr_frac[900] = 10'b0001000100;
    assign isr_frac[901] = 10'b0001000011;
    assign isr_frac[902] = 10'b0001000011;
    assign isr_frac[903] = 10'b0001000010;
    assign isr_frac[904] = 10'b0001000001;
    assign isr_frac[905] = 10'b0001000001;
    assign isr_frac[906] = 10'b0001000000;
    assign isr_frac[907] = 10'b0001000000;
    assign isr_frac[908] = 10'b0000111111;
    assign isr_frac[909] = 10'b0000111110;
    assign isr_frac[910] = 10'b0000111110;
    assign isr_frac[911] = 10'b0000111101;
    assign isr_frac[912] = 10'b0000111101;
    assign isr_frac[913] = 10'b0000111100;
    assign isr_frac[914] = 10'b0000111011;
    assign isr_frac[915] = 10'b0000111011;
    assign isr_frac[916] = 10'b0000111010;
    assign isr_frac[917] = 10'b0000111010;
    assign isr_frac[918] = 10'b0000111001;
    assign isr_frac[919] = 10'b0000111000;
    assign isr_frac[920] = 10'b0000111000;
    assign isr_frac[921] = 10'b0000110111;
    assign isr_frac[922] = 10'b0000110111;
    assign isr_frac[923] = 10'b0000110110;
    assign isr_frac[924] = 10'b0000110101;
    assign isr_frac[925] = 10'b0000110101;
    assign isr_frac[926] = 10'b0000110100;
    assign isr_frac[927] = 10'b0000110100;
    assign isr_frac[928] = 10'b0000110011;
    assign isr_frac[929] = 10'b0000110011;
    assign isr_frac[930] = 10'b0000110010;
    assign isr_frac[931] = 10'b0000110001;
    assign isr_frac[932] = 10'b0000110001;
    assign isr_frac[933] = 10'b0000110000;
    assign isr_frac[934] = 10'b0000110000;
    assign isr_frac[935] = 10'b0000101111;
    assign isr_frac[936] = 10'b0000101111;
    assign isr_frac[937] = 10'b0000101110;
    assign isr_frac[938] = 10'b0000101101;
    assign isr_frac[939] = 10'b0000101101;
    assign isr_frac[940] = 10'b0000101100;
    assign isr_frac[941] = 10'b0000101100;
    assign isr_frac[942] = 10'b0000101011;
    assign isr_frac[943] = 10'b0000101011;
    assign isr_frac[944] = 10'b0000101010;
    assign isr_frac[945] = 10'b0000101001;
    assign isr_frac[946] = 10'b0000101001;
    assign isr_frac[947] = 10'b0000101000;
    assign isr_frac[948] = 10'b0000101000;
    assign isr_frac[949] = 10'b0000100111;
    assign isr_frac[950] = 10'b0000100111;
    assign isr_frac[951] = 10'b0000100110;
    assign isr_frac[952] = 10'b0000100110;
    assign isr_frac[953] = 10'b0000100101;
    assign isr_frac[954] = 10'b0000100100;
    assign isr_frac[955] = 10'b0000100100;
    assign isr_frac[956] = 10'b0000100011;
    assign isr_frac[957] = 10'b0000100011;
    assign isr_frac[958] = 10'b0000100010;
    assign isr_frac[959] = 10'b0000100010;
    assign isr_frac[960] = 10'b0000100001;
    assign isr_frac[961] = 10'b0000100001;
    assign isr_frac[962] = 10'b0000100000;
    assign isr_frac[963] = 10'b0000011111;
    assign isr_frac[964] = 10'b0000011111;
    assign isr_frac[965] = 10'b0000011110;
    assign isr_frac[966] = 10'b0000011110;
    assign isr_frac[967] = 10'b0000011101;
    assign isr_frac[968] = 10'b0000011101;
    assign isr_frac[969] = 10'b0000011100;
    assign isr_frac[970] = 10'b0000011100;
    assign isr_frac[971] = 10'b0000011011;
    assign isr_frac[972] = 10'b0000011011;
    assign isr_frac[973] = 10'b0000011010;
    assign isr_frac[974] = 10'b0000011001;
    assign isr_frac[975] = 10'b0000011001;
    assign isr_frac[976] = 10'b0000011000;
    assign isr_frac[977] = 10'b0000011000;
    assign isr_frac[978] = 10'b0000010111;
    assign isr_frac[979] = 10'b0000010111;
    assign isr_frac[980] = 10'b0000010110;
    assign isr_frac[981] = 10'b0000010110;
    assign isr_frac[982] = 10'b0000010101;
    assign isr_frac[983] = 10'b0000010101;
    assign isr_frac[984] = 10'b0000010100;
    assign isr_frac[985] = 10'b0000010100;
    assign isr_frac[986] = 10'b0000010011;
    assign isr_frac[987] = 10'b0000010011;
    assign isr_frac[988] = 10'b0000010010;
    assign isr_frac[989] = 10'b0000010001;
    assign isr_frac[990] = 10'b0000010001;
    assign isr_frac[991] = 10'b0000010000;
    assign isr_frac[992] = 10'b0000010000;
    assign isr_frac[993] = 10'b0000001111;
    assign isr_frac[994] = 10'b0000001111;
    assign isr_frac[995] = 10'b0000001110;
    assign isr_frac[996] = 10'b0000001110;
    assign isr_frac[997] = 10'b0000001101;
    assign isr_frac[998] = 10'b0000001101;
    assign isr_frac[999] = 10'b0000001100;
    assign isr_frac[1000] = 10'b0000001100;
    assign isr_frac[1001] = 10'b0000001011;
    assign isr_frac[1002] = 10'b0000001011;
    assign isr_frac[1003] = 10'b0000001010;
    assign isr_frac[1004] = 10'b0000001010;
    assign isr_frac[1005] = 10'b0000001001;
    assign isr_frac[1006] = 10'b0000001001;
    assign isr_frac[1007] = 10'b0000001000;
    assign isr_frac[1008] = 10'b0000001000;
    assign isr_frac[1009] = 10'b0000000111;
    assign isr_frac[1010] = 10'b0000000111;
    assign isr_frac[1011] = 10'b0000000110;
    assign isr_frac[1012] = 10'b0000000110;
    assign isr_frac[1013] = 10'b0000000101;
    assign isr_frac[1014] = 10'b0000000101;
    assign isr_frac[1015] = 10'b0000000100;
    assign isr_frac[1016] = 10'b0000000100;
    assign isr_frac[1017] = 10'b0000000011;
    assign isr_frac[1018] = 10'b0000000011;
    assign isr_frac[1019] = 10'b0000000010;
    assign isr_frac[1020] = 10'b0000000010;
    assign isr_frac[1021] = 10'b0000000001;
    assign isr_frac[1022] = 10'b0000000001;
    assign isr_frac[1023] = 10'b0000000000;

assign o_isr = {1'b1, isr_frac[a], 1'b0};// 1.11
assign o_isr_shift_amt = shift_amt[4:1]; // >> 1
assign o_isr_shift_dir = shift_dir;

endmodule