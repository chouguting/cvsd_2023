// list all paths to your design files
`include "../01_RTL/core.v"
`include "../01_RTL/memoryManagementUnit.v"
`include "../01_RTL/indexConverter.v"
`include "../01_RTL/convolutionEngine.v"
`include "../01_RTL/medianFinder.v"
`include "../01_RTL/arctangentApproximator.v"